`define ADDR_BITS 12
`define DATA_BITS 20
`define MUL_DATA_BITS 44
`define SEL_BITS 3
`define KERNAL_NUM 9
`define KERNAL_NUM_1 10
`define KERNAL_NUM_2 11
`define MAX_NUM 3
`define MAX_NUM_1 4
`define IND_BITS 6
`define FALSE 1'b0
`define TRUE 1'b1